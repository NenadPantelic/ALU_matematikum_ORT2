`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:14:01 02/08/2017 
// Design Name: 
// Module Name:    sabiranje 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sabiranje(input [6:0] a,input [6:0] b,output [6:0] z);

assign z = a+b;


endmodule
